--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   14:04:37 01/23/2018
-- Design Name:   
-- Module Name:   C:/Floppy_Bird/Test-Benchs/rng_tb.vhd
-- Project Name:  Floppy_Bird
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: rng
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
USE ieee.numeric_std.ALL;
 
ENTITY rng_tb IS
END rng_tb;
 
ARCHITECTURE behavior OF rng_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT rng
    PORT(
         clk : IN  std_logic;
         rst : IN  std_logic;
         seed : IN  std_logic_vector(9 downto 0);
         random : OUT  std_logic_vector(9 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal clk : std_logic := '0';
   signal rst : std_logic := '0';
   signal seed : std_logic_vector(9 downto 0) := (others => '0');

 	--Outputs
   signal random : std_logic_vector(9 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: rng PORT MAP (
          clk => clk,
          rst => rst,
          seed => seed,
          random => random
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	
		seed <= std_logic_vector(to_unsigned(500,10));
		rst<='1';
      wait for clk_period*10;

      -- insert stimulus here 
		rst <='0';

      wait;
   end process;

END;
